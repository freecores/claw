library verilog;
use verilog.vl_types.all;
entity or1200_wbmux is
    generic(
        width           : integer := 32
    );
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        wb_freeze       : in     vl_logic;
        rfwb_op         : in     vl_logic_vector(2 downto 0);
        rfwb_op2        : in     vl_logic_vector(2 downto 0);
        muxin_a         : in     vl_logic_vector;
        muxin_b         : in     vl_logic_vector;
        muxin_c         : in     vl_logic_vector;
        muxin_d         : in     vl_logic_vector;
        muxin_a2        : in     vl_logic_vector;
        muxin_b2        : in     vl_logic_vector;
        muxin_c2        : in     vl_logic_vector;
        muxin_d2        : in     vl_logic_vector;
        muxout          : out    vl_logic_vector;
        muxreg          : out    vl_logic_vector;
        muxreg_valid    : out    vl_logic;
        muxout2         : out    vl_logic_vector;
        muxreg2         : out    vl_logic_vector;
        muxreg2_valid   : out    vl_logic;
        thread_in       : in     vl_logic_vector(2 downto 0);
        thread_out      : out    vl_logic_vector(2 downto 0)
    );
end or1200_wbmux;

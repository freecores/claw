library verilog;
use verilog.vl_types.all;
entity tb_or1200_rf_top is
    generic(
        aw              : integer := 5;
        dw              : integer := 32
    );
end tb_or1200_rf_top;

library verilog;
use verilog.vl_types.all;
entity tb_or1200_genpc is
end tb_or1200_genpc;

library verilog;
use verilog.vl_types.all;
entity or1200_ctrl is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        id_freeze       : in     vl_logic;
        ex_freeze       : in     vl_logic;
        wb_freeze       : in     vl_logic;
        flushpipe       : in     vl_logic;
        if_insn         : in     vl_logic_vector(31 downto 0);
        ex_insn         : out    vl_logic_vector(31 downto 0);
        branch_op       : out    vl_logic_vector(2 downto 0);
        branch_taken    : in     vl_logic;
        rf_addra        : out    vl_logic_vector(4 downto 0);
        rf_addrb        : out    vl_logic_vector(4 downto 0);
        rf_rda          : out    vl_logic;
        rf_rdb          : out    vl_logic;
        alu_op          : out    vl_logic_vector(3 downto 0);
        mac_op          : out    vl_logic_vector(1 downto 0);
        shrot_op        : out    vl_logic_vector(1 downto 0);
        comp_op         : out    vl_logic_vector(3 downto 0);
        rf_addrw        : out    vl_logic_vector(4 downto 0);
        rfwb_op         : out    vl_logic_vector(2 downto 0);
        wb_insn         : out    vl_logic_vector(31 downto 0);
        simm            : out    vl_logic_vector(31 downto 0);
        branch_addrofs  : out    vl_logic_vector(31 downto 2);
        lsu_addrofs     : out    vl_logic_vector(31 downto 0);
        sel_a           : out    vl_logic_vector(1 downto 0);
        sel_b           : out    vl_logic_vector(1 downto 0);
        lsu_op          : out    vl_logic_vector(3 downto 0);
        cust5_op        : out    vl_logic_vector(4 downto 0);
        cust5_limm      : out    vl_logic_vector(6 downto 0);
        multicycle      : out    vl_logic_vector(1 downto 0);
        spr_addrimm     : out    vl_logic_vector(15 downto 0);
        wbforw_valid    : in     vl_logic;
        du_hwbkpt       : in     vl_logic;
        sig_syscall     : out    vl_logic;
        sig_trap        : out    vl_logic;
        force_dslot_fetch: out    vl_logic;
        no_more_dslot   : out    vl_logic;
        ex_void         : out    vl_logic;
        id_macrc_op     : out    vl_logic;
        ex_macrc_op     : out    vl_logic;
        rfe             : out    vl_logic;
        except_illegal  : out    vl_logic;
        thread_in       : in     vl_logic_vector(2 downto 0);
        thread_out      : out    vl_logic_vector(2 downto 0)
    );
end or1200_ctrl;
